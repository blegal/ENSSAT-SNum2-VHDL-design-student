library IEEE;
use IEEE.std_logic_1164.all;

ENTITY shift_register IS
	PORT ( 
		clock : IN  STD_LOGIC;
		reset : IN  STD_LOGIC;
		load  : IN  STD_LOGIC;
		e     : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		s     : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END shift_register;

ARCHITECTURE behavior OF shift_register IS

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --    

END;