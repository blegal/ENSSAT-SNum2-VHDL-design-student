LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY fonc_logique IS
PORT (
        A : IN  std_logic_vector(3 downto 0);
        B : IN  std_logic_vector(3 downto 0);
        S : OUT std_logic
	);
END fonc_logique;

ARCHITECTURE arch OF fonc_logique IS

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --   

END arch;
