library IEEE;
use IEEE.std_logic_1164.all;

ENTITY led_controler IS 
	PORT ( 
		clock  : IN  STD_LOGIC;
		reset  : IN  STD_LOGIC;
		button : IN  STD_LOGIC;
		red    : OUT STD_LOGIC;
		orange : OUT STD_LOGIC;
		green  : OUT STD_LOGIC
	);
END led_controler;

ARCHITECTURE arch OF led_controler IS

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

END arch;
