library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package conf_counter is

	CONSTANT N    : INTEGER :=   8;
	CONSTANT MINV : INTEGER :=  13;
	CONSTANT MAXV : INTEGER := 222;

end conf_counter;