library IEEE;
use IEEE.std_logic_1164.all;

ENTITY chenillard IS
	PORT ( 
		clock : IN  STD_LOGIC;
		reset : IN  STD_LOGIC;
		s     : OUT STD_LOGIC_VECTOR(7 downto 0)
	);
END chenillard;

ARCHITECTURE behavior OF chenillard IS
    
    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

END;