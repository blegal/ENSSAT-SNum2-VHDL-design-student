LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY logic_alu IS
PORT (
        A : IN  std_logic;
        B : IN  std_logic;
        C : IN  std_logic_vector(2 downto 0);
        D : OUT std_logic
	);
END logic_alu;

ARCHITECTURE arch OF logic_alu IS
BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --   

END arch;
