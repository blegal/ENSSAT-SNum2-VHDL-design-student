LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY adder_4b IS
	PORT (
		A : IN  std_logic_vector(3 downto 0);
		B : IN  std_logic_vector(3 downto 0);
		S : OUT std_logic_vector(4 downto 0)
	);
END adder_4b;

ARCHITECTURE arch OF adder_4b IS


    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --
    

BEGIN

    --
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    -- ... ... ... ... ... ...
    --

END arch;
